-- trolley_system.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity trolley_system is
	port (
		altpll_0_c1_clk                          : out   std_logic;                                        --                       altpll_0_c1.clk
		button_button_external_connection_export : in    std_logic                     := '0';             -- button_button_external_connection.export
		button_led_external_connection_export    : out   std_logic;                                        --    button_led_external_connection.export
		cam_uart_external_connection_rxd         : in    std_logic                     := '0';             --      cam_uart_external_connection.rxd
		cam_uart_external_connection_txd         : out   std_logic;                                        --                                  .txd
		clk_clk                                  : in    std_logic                     := '0';             --                               clk.clk
		epcs_flash_controller_0_external_dclk    : out   std_logic;                                        --  epcs_flash_controller_0_external.dclk
		epcs_flash_controller_0_external_sce     : out   std_logic;                                        --                                  .sce
		epcs_flash_controller_0_external_sdo     : out   std_logic;                                        --                                  .sdo
		epcs_flash_controller_0_external_data0   : in    std_logic                     := '0';             --                                  .data0
		green_leds_external_connection_export    : out   std_logic_vector(7 downto 0);                     --    green_leds_external_connection.export
		key_external_connection_export           : in    std_logic                     := '0';             --           key_external_connection.export
		motor_l_external_connection_export       : out   std_logic_vector(2 downto 0);                     --       motor_l_external_connection.export
		motor_r_external_connection_export       : out   std_logic_vector(2 downto 0);                     --       motor_r_external_connection.export
		prox_sensor_external_connection_export   : in    std_logic                     := '0';             --   prox_sensor_external_connection.export
		reset_reset_n                            : in    std_logic                     := '0';             --                             reset.reset_n
		sdram_controller_0_wire_addr             : out   std_logic_vector(11 downto 0);                    --           sdram_controller_0_wire.addr
		sdram_controller_0_wire_ba               : out   std_logic_vector(1 downto 0);                     --                                  .ba
		sdram_controller_0_wire_cas_n            : out   std_logic;                                        --                                  .cas_n
		sdram_controller_0_wire_cke              : out   std_logic;                                        --                                  .cke
		sdram_controller_0_wire_cs_n             : out   std_logic;                                        --                                  .cs_n
		sdram_controller_0_wire_dq               : inout std_logic_vector(15 downto 0) := (others => '0'); --                                  .dq
		sdram_controller_0_wire_dqm              : out   std_logic_vector(1 downto 0);                     --                                  .dqm
		sdram_controller_0_wire_ras_n            : out   std_logic;                                        --                                  .ras_n
		sdram_controller_0_wire_we_n             : out   std_logic;                                        --                                  .we_n
		speaker_external_connection_export       : out   std_logic;                                        --       speaker_external_connection.export
		wifi_uart_external_connection_rxd        : in    std_logic                     := '0';             --     wifi_uart_external_connection.rxd
		wifi_uart_external_connection_txd        : out   std_logic                                         --                                  .txd
	);
end entity trolley_system;

architecture rtl of trolley_system is
	component trolley_system_altpll_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component trolley_system_altpll_0;

	component trolley_system_button_button is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component trolley_system_button_button;

	component trolley_system_button_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component trolley_system_button_led;

	component trolley_system_cam_uart is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component trolley_system_cam_uart;

	component trolley_system_epcs_flash_controller_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			address    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read_n     : in  std_logic                     := 'X';             -- read_n
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			irq        : out std_logic;                                        -- irq
			dclk       : out std_logic;                                        -- export
			sce        : out std_logic;                                        -- export
			sdo        : out std_logic;                                        -- export
			data0      : in  std_logic                     := 'X'              -- export
		);
	end component trolley_system_epcs_flash_controller_0;

	component trolley_system_green_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component trolley_system_green_leds;

	component trolley_system_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component trolley_system_jtag_uart_0;

	component trolley_system_motor_l is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(2 downto 0)                      -- export
		);
	end component trolley_system_motor_l;

	component trolley_system_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(24 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(24 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component trolley_system_nios2_gen2_0;

	component trolley_system_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component trolley_system_onchip_memory2_0;

	component trolley_system_sdram_controller_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component trolley_system_sdram_controller_0;

	component trolley_system_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component trolley_system_sysid_qsys_0;

	component trolley_system_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component trolley_system_timer_0;

	component trolley_system_wifi_uart is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component trolley_system_wifi_uart;

	component trolley_system_mm_interconnect_0 is
		port (
			altpll_0_c0_clk                                      : in  std_logic                     := 'X';             -- clk
			key_reset_reset_bridge_in_reset_reset                : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                     : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                 : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                        : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                    : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                       : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                 : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest          : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                 : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			button_button_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			button_button_s1_write                               : out std_logic;                                        -- write
			button_button_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			button_button_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			button_button_s1_chipselect                          : out std_logic;                                        -- chipselect
			button_led_s1_address                                : out std_logic_vector(1 downto 0);                     -- address
			button_led_s1_write                                  : out std_logic;                                        -- write
			button_led_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			button_led_s1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			button_led_s1_chipselect                             : out std_logic;                                        -- chipselect
			cam_uart_s1_address                                  : out std_logic_vector(2 downto 0);                     -- address
			cam_uart_s1_write                                    : out std_logic;                                        -- write
			cam_uart_s1_read                                     : out std_logic;                                        -- read
			cam_uart_s1_readdata                                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			cam_uart_s1_writedata                                : out std_logic_vector(15 downto 0);                    -- writedata
			cam_uart_s1_begintransfer                            : out std_logic;                                        -- begintransfer
			cam_uart_s1_chipselect                               : out std_logic;                                        -- chipselect
			epcs_flash_controller_0_epcs_control_port_address    : out std_logic_vector(8 downto 0);                     -- address
			epcs_flash_controller_0_epcs_control_port_write      : out std_logic;                                        -- write
			epcs_flash_controller_0_epcs_control_port_read       : out std_logic;                                        -- read
			epcs_flash_controller_0_epcs_control_port_readdata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			epcs_flash_controller_0_epcs_control_port_writedata  : out std_logic_vector(31 downto 0);                    -- writedata
			epcs_flash_controller_0_epcs_control_port_chipselect : out std_logic;                                        -- chipselect
			green_leds_s1_address                                : out std_logic_vector(1 downto 0);                     -- address
			green_leds_s1_write                                  : out std_logic;                                        -- write
			green_leds_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			green_leds_s1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			green_leds_s1_chipselect                             : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address                : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                  : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                   : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect             : out std_logic;                                        -- chipselect
			key_s1_address                                       : out std_logic_vector(1 downto 0);                     -- address
			key_s1_write                                         : out std_logic;                                        -- write
			key_s1_readdata                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			key_s1_writedata                                     : out std_logic_vector(31 downto 0);                    -- writedata
			key_s1_chipselect                                    : out std_logic;                                        -- chipselect
			motor_l_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			motor_l_s1_write                                     : out std_logic;                                        -- write
			motor_l_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			motor_l_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			motor_l_s1_chipselect                                : out std_logic;                                        -- chipselect
			motor_r_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			motor_r_s1_write                                     : out std_logic;                                        -- write
			motor_r_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			motor_r_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			motor_r_s1_chipselect                                : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address                 : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                   : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                    : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable              : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest             : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess             : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                          : out std_logic_vector(11 downto 0);                    -- address
			onchip_memory2_0_s1_write                            : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                       : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                            : out std_logic;                                        -- clken
			prox_sensor_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			prox_sensor_s1_write                                 : out std_logic;                                        -- write
			prox_sensor_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			prox_sensor_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			prox_sensor_s1_chipselect                            : out std_logic;                                        -- chipselect
			sdram_controller_0_s1_address                        : out std_logic_vector(21 downto 0);                    -- address
			sdram_controller_0_s1_write                          : out std_logic;                                        -- write
			sdram_controller_0_s1_read                           : out std_logic;                                        -- read
			sdram_controller_0_s1_readdata                       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_controller_0_s1_writedata                      : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_controller_0_s1_byteenable                     : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_controller_0_s1_readdatavalid                  : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_0_s1_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_0_s1_chipselect                     : out std_logic;                                        -- chipselect
			speaker_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			speaker_s1_write                                     : out std_logic;                                        -- write
			speaker_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			speaker_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			speaker_s1_chipselect                                : out std_logic;                                        -- chipselect
			sysid_qsys_0_control_slave_address                   : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                                   : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                     : out std_logic;                                        -- write
			timer_0_s1_readdata                                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                                 : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                                : out std_logic;                                        -- chipselect
			wifi_uart_s1_address                                 : out std_logic_vector(2 downto 0);                     -- address
			wifi_uart_s1_write                                   : out std_logic;                                        -- write
			wifi_uart_s1_read                                    : out std_logic;                                        -- read
			wifi_uart_s1_readdata                                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			wifi_uart_s1_writedata                               : out std_logic_vector(15 downto 0);                    -- writedata
			wifi_uart_s1_begintransfer                           : out std_logic;                                        -- begintransfer
			wifi_uart_s1_chipselect                              : out std_logic                                         -- chipselect
		);
	end component trolley_system_mm_interconnect_0;

	component trolley_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			receiver6_irq : in  std_logic                     := 'X'; -- irq
			receiver7_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component trolley_system_irq_mapper;

	component trolley_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component trolley_system_rst_controller;

	component trolley_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component trolley_system_rst_controller_001;

	component trolley_system_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component trolley_system_rst_controller_002;

	signal altpll_0_c0_clk                                                             : std_logic;                     -- altpll_0:c0 -> [button_button:clk, button_led:clk, cam_uart:clk, epcs_flash_controller_0:clk, green_leds:clk, irq_mapper:clk, jtag_uart_0:clk, key:clk, mm_interconnect_0:altpll_0_c0_clk, motor_l:clk, motor_r:clk, nios2_gen2_0:clk, onchip_memory2_0:clk, prox_sensor:clk, rst_controller_001:clk, rst_controller_002:clk, sdram_controller_0:clk, speaker:clk, sysid_qsys_0:clock, timer_0:clk, wifi_uart:clk]
	signal nios2_gen2_0_data_master_readdata                                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                        : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                        : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                            : std_logic_vector(24 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                         : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                               : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                              : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                          : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                                 : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                                     : std_logic_vector(24 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                        : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect                  : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata                    : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest                 : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address                     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read                        : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write                       : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata                       : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address                        : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata                     : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest                  : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess                  : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address                      : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read                         : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable                   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write                        : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_chipselect      : std_logic;                     -- mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_chipselect -> epcs_flash_controller_0:chipselect
	signal mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_readdata        : std_logic_vector(31 downto 0); -- epcs_flash_controller_0:readdata -> mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_readdata
	signal mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_address         : std_logic_vector(8 downto 0);  -- mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_address -> epcs_flash_controller_0:address
	signal mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read            : std_logic;                     -- mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_read -> mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read:in
	signal mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write           : std_logic;                     -- mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_write -> mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write:in
	signal mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_writedata -> epcs_flash_controller_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                              : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                               : std_logic_vector(11 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                                 : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                                 : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_sdram_controller_0_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_chipselect -> sdram_controller_0:az_cs
	signal mm_interconnect_0_sdram_controller_0_s1_readdata                            : std_logic_vector(15 downto 0); -- sdram_controller_0:za_data -> mm_interconnect_0:sdram_controller_0_s1_readdata
	signal mm_interconnect_0_sdram_controller_0_s1_waitrequest                         : std_logic;                     -- sdram_controller_0:za_waitrequest -> mm_interconnect_0:sdram_controller_0_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_0_s1_address                             : std_logic_vector(21 downto 0); -- mm_interconnect_0:sdram_controller_0_s1_address -> sdram_controller_0:az_addr
	signal mm_interconnect_0_sdram_controller_0_s1_read                                : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_read -> mm_interconnect_0_sdram_controller_0_s1_read:in
	signal mm_interconnect_0_sdram_controller_0_s1_byteenable                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_controller_0_s1_byteenable -> mm_interconnect_0_sdram_controller_0_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_0_s1_readdatavalid                       : std_logic;                     -- sdram_controller_0:za_valid -> mm_interconnect_0:sdram_controller_0_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_0_s1_write                               : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_write -> mm_interconnect_0_sdram_controller_0_s1_write:in
	signal mm_interconnect_0_sdram_controller_0_s1_writedata                           : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_controller_0_s1_writedata -> sdram_controller_0:az_data
	signal mm_interconnect_0_cam_uart_s1_chipselect                                    : std_logic;                     -- mm_interconnect_0:cam_uart_s1_chipselect -> cam_uart:chipselect
	signal mm_interconnect_0_cam_uart_s1_readdata                                      : std_logic_vector(15 downto 0); -- cam_uart:readdata -> mm_interconnect_0:cam_uart_s1_readdata
	signal mm_interconnect_0_cam_uart_s1_address                                       : std_logic_vector(2 downto 0);  -- mm_interconnect_0:cam_uart_s1_address -> cam_uart:address
	signal mm_interconnect_0_cam_uart_s1_read                                          : std_logic;                     -- mm_interconnect_0:cam_uart_s1_read -> mm_interconnect_0_cam_uart_s1_read:in
	signal mm_interconnect_0_cam_uart_s1_begintransfer                                 : std_logic;                     -- mm_interconnect_0:cam_uart_s1_begintransfer -> cam_uart:begintransfer
	signal mm_interconnect_0_cam_uart_s1_write                                         : std_logic;                     -- mm_interconnect_0:cam_uart_s1_write -> mm_interconnect_0_cam_uart_s1_write:in
	signal mm_interconnect_0_cam_uart_s1_writedata                                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:cam_uart_s1_writedata -> cam_uart:writedata
	signal mm_interconnect_0_wifi_uart_s1_chipselect                                   : std_logic;                     -- mm_interconnect_0:wifi_uart_s1_chipselect -> wifi_uart:chipselect
	signal mm_interconnect_0_wifi_uart_s1_readdata                                     : std_logic_vector(15 downto 0); -- wifi_uart:readdata -> mm_interconnect_0:wifi_uart_s1_readdata
	signal mm_interconnect_0_wifi_uart_s1_address                                      : std_logic_vector(2 downto 0);  -- mm_interconnect_0:wifi_uart_s1_address -> wifi_uart:address
	signal mm_interconnect_0_wifi_uart_s1_read                                         : std_logic;                     -- mm_interconnect_0:wifi_uart_s1_read -> mm_interconnect_0_wifi_uart_s1_read:in
	signal mm_interconnect_0_wifi_uart_s1_begintransfer                                : std_logic;                     -- mm_interconnect_0:wifi_uart_s1_begintransfer -> wifi_uart:begintransfer
	signal mm_interconnect_0_wifi_uart_s1_write                                        : std_logic;                     -- mm_interconnect_0:wifi_uart_s1_write -> mm_interconnect_0_wifi_uart_s1_write:in
	signal mm_interconnect_0_wifi_uart_s1_writedata                                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:wifi_uart_s1_writedata -> wifi_uart:writedata
	signal mm_interconnect_0_prox_sensor_s1_chipselect                                 : std_logic;                     -- mm_interconnect_0:prox_sensor_s1_chipselect -> prox_sensor:chipselect
	signal mm_interconnect_0_prox_sensor_s1_readdata                                   : std_logic_vector(31 downto 0); -- prox_sensor:readdata -> mm_interconnect_0:prox_sensor_s1_readdata
	signal mm_interconnect_0_prox_sensor_s1_address                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:prox_sensor_s1_address -> prox_sensor:address
	signal mm_interconnect_0_prox_sensor_s1_write                                      : std_logic;                     -- mm_interconnect_0:prox_sensor_s1_write -> mm_interconnect_0_prox_sensor_s1_write:in
	signal mm_interconnect_0_prox_sensor_s1_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:prox_sensor_s1_writedata -> prox_sensor:writedata
	signal mm_interconnect_0_motor_r_s1_chipselect                                     : std_logic;                     -- mm_interconnect_0:motor_r_s1_chipselect -> motor_r:chipselect
	signal mm_interconnect_0_motor_r_s1_readdata                                       : std_logic_vector(31 downto 0); -- motor_r:readdata -> mm_interconnect_0:motor_r_s1_readdata
	signal mm_interconnect_0_motor_r_s1_address                                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:motor_r_s1_address -> motor_r:address
	signal mm_interconnect_0_motor_r_s1_write                                          : std_logic;                     -- mm_interconnect_0:motor_r_s1_write -> mm_interconnect_0_motor_r_s1_write:in
	signal mm_interconnect_0_motor_r_s1_writedata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:motor_r_s1_writedata -> motor_r:writedata
	signal mm_interconnect_0_motor_l_s1_chipselect                                     : std_logic;                     -- mm_interconnect_0:motor_l_s1_chipselect -> motor_l:chipselect
	signal mm_interconnect_0_motor_l_s1_readdata                                       : std_logic_vector(31 downto 0); -- motor_l:readdata -> mm_interconnect_0:motor_l_s1_readdata
	signal mm_interconnect_0_motor_l_s1_address                                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:motor_l_s1_address -> motor_l:address
	signal mm_interconnect_0_motor_l_s1_write                                          : std_logic;                     -- mm_interconnect_0:motor_l_s1_write -> mm_interconnect_0_motor_l_s1_write:in
	signal mm_interconnect_0_motor_l_s1_writedata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:motor_l_s1_writedata -> motor_l:writedata
	signal mm_interconnect_0_green_leds_s1_chipselect                                  : std_logic;                     -- mm_interconnect_0:green_leds_s1_chipselect -> green_leds:chipselect
	signal mm_interconnect_0_green_leds_s1_readdata                                    : std_logic_vector(31 downto 0); -- green_leds:readdata -> mm_interconnect_0:green_leds_s1_readdata
	signal mm_interconnect_0_green_leds_s1_address                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:green_leds_s1_address -> green_leds:address
	signal mm_interconnect_0_green_leds_s1_write                                       : std_logic;                     -- mm_interconnect_0:green_leds_s1_write -> mm_interconnect_0_green_leds_s1_write:in
	signal mm_interconnect_0_green_leds_s1_writedata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:green_leds_s1_writedata -> green_leds:writedata
	signal mm_interconnect_0_button_button_s1_chipselect                               : std_logic;                     -- mm_interconnect_0:button_button_s1_chipselect -> button_button:chipselect
	signal mm_interconnect_0_button_button_s1_readdata                                 : std_logic_vector(31 downto 0); -- button_button:readdata -> mm_interconnect_0:button_button_s1_readdata
	signal mm_interconnect_0_button_button_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:button_button_s1_address -> button_button:address
	signal mm_interconnect_0_button_button_s1_write                                    : std_logic;                     -- mm_interconnect_0:button_button_s1_write -> mm_interconnect_0_button_button_s1_write:in
	signal mm_interconnect_0_button_button_s1_writedata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:button_button_s1_writedata -> button_button:writedata
	signal mm_interconnect_0_button_led_s1_chipselect                                  : std_logic;                     -- mm_interconnect_0:button_led_s1_chipselect -> button_led:chipselect
	signal mm_interconnect_0_button_led_s1_readdata                                    : std_logic_vector(31 downto 0); -- button_led:readdata -> mm_interconnect_0:button_led_s1_readdata
	signal mm_interconnect_0_button_led_s1_address                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:button_led_s1_address -> button_led:address
	signal mm_interconnect_0_button_led_s1_write                                       : std_logic;                     -- mm_interconnect_0:button_led_s1_write -> mm_interconnect_0_button_led_s1_write:in
	signal mm_interconnect_0_button_led_s1_writedata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:button_led_s1_writedata -> button_led:writedata
	signal mm_interconnect_0_speaker_s1_chipselect                                     : std_logic;                     -- mm_interconnect_0:speaker_s1_chipselect -> speaker:chipselect
	signal mm_interconnect_0_speaker_s1_readdata                                       : std_logic_vector(31 downto 0); -- speaker:readdata -> mm_interconnect_0:speaker_s1_readdata
	signal mm_interconnect_0_speaker_s1_address                                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:speaker_s1_address -> speaker:address
	signal mm_interconnect_0_speaker_s1_write                                          : std_logic;                     -- mm_interconnect_0:speaker_s1_write -> mm_interconnect_0_speaker_s1_write:in
	signal mm_interconnect_0_speaker_s1_writedata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:speaker_s1_writedata -> speaker:writedata
	signal mm_interconnect_0_timer_0_s1_chipselect                                     : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                                       : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                                          : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_key_s1_chipselect                                         : std_logic;                     -- mm_interconnect_0:key_s1_chipselect -> key:chipselect
	signal mm_interconnect_0_key_s1_readdata                                           : std_logic_vector(31 downto 0); -- key:readdata -> mm_interconnect_0:key_s1_readdata
	signal mm_interconnect_0_key_s1_address                                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:key_s1_address -> key:address
	signal mm_interconnect_0_key_s1_write                                              : std_logic;                     -- mm_interconnect_0:key_s1_write -> mm_interconnect_0_key_s1_write:in
	signal mm_interconnect_0_key_s1_writedata                                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:key_s1_writedata -> key:writedata
	signal irq_mapper_receiver0_irq                                                    : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                    : std_logic;                     -- cam_uart:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                    : std_logic;                     -- wifi_uart:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                    : std_logic;                     -- prox_sensor:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                                    : std_logic;                     -- button_button:irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                                    : std_logic;                     -- timer_0:irq -> irq_mapper:receiver5_irq
	signal irq_mapper_receiver6_irq                                                    : std_logic;                     -- epcs_flash_controller_0:irq -> irq_mapper:receiver6_irq
	signal irq_mapper_receiver7_irq                                                    : std_logic;                     -- key:irq -> irq_mapper:receiver7_irq
	signal nios2_gen2_0_irq_irq                                                        : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                              : std_logic;                     -- rst_controller:reset_out -> altpll_0:reset
	signal nios2_gen2_0_debug_reset_request_reset                                      : std_logic;                     -- nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                                          : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_001_reset_out_reset_req                                      : std_logic;                     -- rst_controller_001:reset_req -> [epcs_flash_controller_0:reset_req, nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal rst_controller_002_reset_out_reset                                          : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:key_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                                     : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv              : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv             : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read_ports_inv  : std_logic;                     -- mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read:inv -> epcs_flash_controller_0:read_n
	signal mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write_ports_inv : std_logic;                     -- mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write:inv -> epcs_flash_controller_0:write_n
	signal mm_interconnect_0_sdram_controller_0_s1_read_ports_inv                      : std_logic;                     -- mm_interconnect_0_sdram_controller_0_s1_read:inv -> sdram_controller_0:az_rd_n
	signal mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv                : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_controller_0_s1_byteenable:inv -> sdram_controller_0:az_be_n
	signal mm_interconnect_0_sdram_controller_0_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_sdram_controller_0_s1_write:inv -> sdram_controller_0:az_wr_n
	signal mm_interconnect_0_cam_uart_s1_read_ports_inv                                : std_logic;                     -- mm_interconnect_0_cam_uart_s1_read:inv -> cam_uart:read_n
	signal mm_interconnect_0_cam_uart_s1_write_ports_inv                               : std_logic;                     -- mm_interconnect_0_cam_uart_s1_write:inv -> cam_uart:write_n
	signal mm_interconnect_0_wifi_uart_s1_read_ports_inv                               : std_logic;                     -- mm_interconnect_0_wifi_uart_s1_read:inv -> wifi_uart:read_n
	signal mm_interconnect_0_wifi_uart_s1_write_ports_inv                              : std_logic;                     -- mm_interconnect_0_wifi_uart_s1_write:inv -> wifi_uart:write_n
	signal mm_interconnect_0_prox_sensor_s1_write_ports_inv                            : std_logic;                     -- mm_interconnect_0_prox_sensor_s1_write:inv -> prox_sensor:write_n
	signal mm_interconnect_0_motor_r_s1_write_ports_inv                                : std_logic;                     -- mm_interconnect_0_motor_r_s1_write:inv -> motor_r:write_n
	signal mm_interconnect_0_motor_l_s1_write_ports_inv                                : std_logic;                     -- mm_interconnect_0_motor_l_s1_write:inv -> motor_l:write_n
	signal mm_interconnect_0_green_leds_s1_write_ports_inv                             : std_logic;                     -- mm_interconnect_0_green_leds_s1_write:inv -> green_leds:write_n
	signal mm_interconnect_0_button_button_s1_write_ports_inv                          : std_logic;                     -- mm_interconnect_0_button_button_s1_write:inv -> button_button:write_n
	signal mm_interconnect_0_button_led_s1_write_ports_inv                             : std_logic;                     -- mm_interconnect_0_button_led_s1_write:inv -> button_led:write_n
	signal mm_interconnect_0_speaker_s1_write_ports_inv                                : std_logic;                     -- mm_interconnect_0_speaker_s1_write:inv -> speaker:write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                                : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_key_s1_write_ports_inv                                    : std_logic;                     -- mm_interconnect_0_key_s1_write:inv -> key:write_n
	signal rst_controller_001_reset_out_reset_ports_inv                                : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [button_button:reset_n, button_led:reset_n, cam_uart:reset_n, epcs_flash_controller_0:reset_n, green_leds:reset_n, jtag_uart_0:rst_n, motor_l:reset_n, motor_r:reset_n, nios2_gen2_0:reset_n, prox_sensor:reset_n, sdram_controller_0:reset_n, speaker:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n, wifi_uart:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                                : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> key:reset_n

begin

	altpll_0 : component trolley_system_altpll_0
		port map (
			clk                => clk_clk,                        --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset, -- inclk_interface_reset.reset
			read               => open,                           --             pll_slave.read
			write              => open,                           --                      .write
			address            => open,                           --                      .address
			readdata           => open,                           --                      .readdata
			writedata          => open,                           --                      .writedata
			c0                 => altpll_0_c0_clk,                --                    c0.clk
			c1                 => altpll_0_c1_clk,                --                    c1.clk
			scandone           => open,                           --           (terminated)
			scandataout        => open,                           --           (terminated)
			areset             => '0',                            --           (terminated)
			locked             => open,                           --           (terminated)
			phasedone          => open,                           --           (terminated)
			phasecounterselect => "0000",                         --           (terminated)
			phaseupdown        => '0',                            --           (terminated)
			phasestep          => '0',                            --           (terminated)
			scanclk            => '0',                            --           (terminated)
			scanclkena         => '0',                            --           (terminated)
			scandata           => '0',                            --           (terminated)
			configupdate       => '0'                             --           (terminated)
		);

	button_button : component trolley_system_button_button
		port map (
			clk        => altpll_0_c0_clk,                                    --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_button_button_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_button_button_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_button_button_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_button_button_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_button_button_s1_readdata,        --                    .readdata
			in_port    => button_button_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver4_irq                            --                 irq.irq
		);

	button_led : component trolley_system_button_led
		port map (
			clk        => altpll_0_c0_clk,                                 --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_button_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_button_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_button_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_button_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_button_led_s1_readdata,        --                    .readdata
			out_port   => button_led_external_connection_export            -- external_connection.export
		);

	cam_uart : component trolley_system_cam_uart
		port map (
			clk           => altpll_0_c0_clk,                               --                 clk.clk
			reset_n       => rst_controller_001_reset_out_reset_ports_inv,  --               reset.reset_n
			address       => mm_interconnect_0_cam_uart_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_cam_uart_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_cam_uart_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_cam_uart_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_cam_uart_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_cam_uart_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_cam_uart_s1_readdata,        --                    .readdata
			rxd           => cam_uart_external_connection_rxd,              -- external_connection.export
			txd           => cam_uart_external_connection_txd,              --                    .export
			irq           => irq_mapper_receiver1_irq                       --                 irq.irq
		);

	epcs_flash_controller_0 : component trolley_system_epcs_flash_controller_0
		port map (
			clk        => altpll_0_c0_clk,                                                             --               clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,                                --             reset.reset_n
			reset_req  => rst_controller_001_reset_out_reset_req,                                      --                  .reset_req
			address    => mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_address,         -- epcs_control_port.address
			chipselect => mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_chipselect,      --                  .chipselect
			read_n     => mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read_ports_inv,  --                  .read_n
			readdata   => mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_readdata,        --                  .readdata
			write_n    => mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write_ports_inv, --                  .write_n
			writedata  => mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_writedata,       --                  .writedata
			irq        => irq_mapper_receiver6_irq,                                                    --               irq.irq
			dclk       => epcs_flash_controller_0_external_dclk,                                       --          external.export
			sce        => epcs_flash_controller_0_external_sce,                                        --                  .export
			sdo        => epcs_flash_controller_0_external_sdo,                                        --                  .export
			data0      => epcs_flash_controller_0_external_data0                                       --                  .export
		);

	green_leds : component trolley_system_green_leds
		port map (
			clk        => altpll_0_c0_clk,                                 --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_green_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_green_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_green_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_green_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_green_leds_s1_readdata,        --                    .readdata
			out_port   => green_leds_external_connection_export            -- external_connection.export
		);

	jtag_uart_0 : component trolley_system_jtag_uart_0
		port map (
			clk            => altpll_0_c0_clk,                                                 --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	key : component trolley_system_button_button
		port map (
			clk        => altpll_0_c0_clk,                              --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_key_s1_address,             --                  s1.address
			write_n    => mm_interconnect_0_key_s1_write_ports_inv,     --                    .write_n
			writedata  => mm_interconnect_0_key_s1_writedata,           --                    .writedata
			chipselect => mm_interconnect_0_key_s1_chipselect,          --                    .chipselect
			readdata   => mm_interconnect_0_key_s1_readdata,            --                    .readdata
			in_port    => key_external_connection_export,               -- external_connection.export
			irq        => irq_mapper_receiver7_irq                      --                 irq.irq
		);

	motor_l : component trolley_system_motor_l
		port map (
			clk        => altpll_0_c0_clk,                              --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_motor_l_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_motor_l_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_motor_l_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_motor_l_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_motor_l_s1_readdata,        --                    .readdata
			out_port   => motor_l_external_connection_export            -- external_connection.export
		);

	motor_r : component trolley_system_motor_l
		port map (
			clk        => altpll_0_c0_clk,                              --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_motor_r_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_motor_r_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_motor_r_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_motor_r_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_motor_r_s1_readdata,        --                    .readdata
			out_port   => motor_r_external_connection_export            -- external_connection.export
		);

	nios2_gen2_0 : component trolley_system_nios2_gen2_0
		port map (
			clk                                 => altpll_0_c0_clk,                                            --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,               --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,                     --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component trolley_system_onchip_memory2_0
		port map (
			clk        => altpll_0_c0_clk,                                  --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,               -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req,           --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	prox_sensor : component trolley_system_button_button
		port map (
			clk        => altpll_0_c0_clk,                                  --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_prox_sensor_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_prox_sensor_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_prox_sensor_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_prox_sensor_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_prox_sensor_s1_readdata,        --                    .readdata
			in_port    => prox_sensor_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver3_irq                          --                 irq.irq
		);

	sdram_controller_0 : component trolley_system_sdram_controller_0
		port map (
			clk            => altpll_0_c0_clk,                                              --   clk.clk
			reset_n        => rst_controller_001_reset_out_reset_ports_inv,                 -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_0_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_0_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_0_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_0_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_0_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_0_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_0_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_0_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_controller_0_wire_addr,                                 --  wire.export
			zs_ba          => sdram_controller_0_wire_ba,                                   --      .export
			zs_cas_n       => sdram_controller_0_wire_cas_n,                                --      .export
			zs_cke         => sdram_controller_0_wire_cke,                                  --      .export
			zs_cs_n        => sdram_controller_0_wire_cs_n,                                 --      .export
			zs_dq          => sdram_controller_0_wire_dq,                                   --      .export
			zs_dqm         => sdram_controller_0_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_controller_0_wire_ras_n,                                --      .export
			zs_we_n        => sdram_controller_0_wire_we_n                                  --      .export
		);

	speaker : component trolley_system_button_led
		port map (
			clk        => altpll_0_c0_clk,                              --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_speaker_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_speaker_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_speaker_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_speaker_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_speaker_s1_readdata,        --                    .readdata
			out_port   => speaker_external_connection_export            -- external_connection.export
		);

	sysid_qsys_0 : component trolley_system_sysid_qsys_0
		port map (
			clock    => altpll_0_c0_clk,                                         --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,            --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	timer_0 : component trolley_system_timer_0
		port map (
			clk        => altpll_0_c0_clk,                              --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver5_irq                      --   irq.irq
		);

	wifi_uart : component trolley_system_wifi_uart
		port map (
			clk           => altpll_0_c0_clk,                                --                 clk.clk
			reset_n       => rst_controller_001_reset_out_reset_ports_inv,   --               reset.reset_n
			address       => mm_interconnect_0_wifi_uart_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_wifi_uart_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_wifi_uart_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_wifi_uart_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_wifi_uart_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_wifi_uart_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_wifi_uart_s1_readdata,        --                    .readdata
			rxd           => wifi_uart_external_connection_rxd,              -- external_connection.export
			txd           => wifi_uart_external_connection_txd,              --                    .export
			irq           => irq_mapper_receiver2_irq                        --                 irq.irq
		);

	mm_interconnect_0 : component trolley_system_mm_interconnect_0
		port map (
			altpll_0_c0_clk                                      => altpll_0_c0_clk,                                                        --                               altpll_0_c0.clk
			key_reset_reset_bridge_in_reset_reset                => rst_controller_002_reset_out_reset,                                     --           key_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset       => rst_controller_001_reset_out_reset,                                     --  nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                     => nios2_gen2_0_data_master_address,                                       --                  nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                 => nios2_gen2_0_data_master_waitrequest,                                   --                                          .waitrequest
			nios2_gen2_0_data_master_byteenable                  => nios2_gen2_0_data_master_byteenable,                                    --                                          .byteenable
			nios2_gen2_0_data_master_read                        => nios2_gen2_0_data_master_read,                                          --                                          .read
			nios2_gen2_0_data_master_readdata                    => nios2_gen2_0_data_master_readdata,                                      --                                          .readdata
			nios2_gen2_0_data_master_write                       => nios2_gen2_0_data_master_write,                                         --                                          .write
			nios2_gen2_0_data_master_writedata                   => nios2_gen2_0_data_master_writedata,                                     --                                          .writedata
			nios2_gen2_0_data_master_debugaccess                 => nios2_gen2_0_data_master_debugaccess,                                   --                                          .debugaccess
			nios2_gen2_0_instruction_master_address              => nios2_gen2_0_instruction_master_address,                                --           nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest          => nios2_gen2_0_instruction_master_waitrequest,                            --                                          .waitrequest
			nios2_gen2_0_instruction_master_read                 => nios2_gen2_0_instruction_master_read,                                   --                                          .read
			nios2_gen2_0_instruction_master_readdata             => nios2_gen2_0_instruction_master_readdata,                               --                                          .readdata
			button_button_s1_address                             => mm_interconnect_0_button_button_s1_address,                             --                          button_button_s1.address
			button_button_s1_write                               => mm_interconnect_0_button_button_s1_write,                               --                                          .write
			button_button_s1_readdata                            => mm_interconnect_0_button_button_s1_readdata,                            --                                          .readdata
			button_button_s1_writedata                           => mm_interconnect_0_button_button_s1_writedata,                           --                                          .writedata
			button_button_s1_chipselect                          => mm_interconnect_0_button_button_s1_chipselect,                          --                                          .chipselect
			button_led_s1_address                                => mm_interconnect_0_button_led_s1_address,                                --                             button_led_s1.address
			button_led_s1_write                                  => mm_interconnect_0_button_led_s1_write,                                  --                                          .write
			button_led_s1_readdata                               => mm_interconnect_0_button_led_s1_readdata,                               --                                          .readdata
			button_led_s1_writedata                              => mm_interconnect_0_button_led_s1_writedata,                              --                                          .writedata
			button_led_s1_chipselect                             => mm_interconnect_0_button_led_s1_chipselect,                             --                                          .chipselect
			cam_uart_s1_address                                  => mm_interconnect_0_cam_uart_s1_address,                                  --                               cam_uart_s1.address
			cam_uart_s1_write                                    => mm_interconnect_0_cam_uart_s1_write,                                    --                                          .write
			cam_uart_s1_read                                     => mm_interconnect_0_cam_uart_s1_read,                                     --                                          .read
			cam_uart_s1_readdata                                 => mm_interconnect_0_cam_uart_s1_readdata,                                 --                                          .readdata
			cam_uart_s1_writedata                                => mm_interconnect_0_cam_uart_s1_writedata,                                --                                          .writedata
			cam_uart_s1_begintransfer                            => mm_interconnect_0_cam_uart_s1_begintransfer,                            --                                          .begintransfer
			cam_uart_s1_chipselect                               => mm_interconnect_0_cam_uart_s1_chipselect,                               --                                          .chipselect
			epcs_flash_controller_0_epcs_control_port_address    => mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_address,    -- epcs_flash_controller_0_epcs_control_port.address
			epcs_flash_controller_0_epcs_control_port_write      => mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write,      --                                          .write
			epcs_flash_controller_0_epcs_control_port_read       => mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read,       --                                          .read
			epcs_flash_controller_0_epcs_control_port_readdata   => mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_readdata,   --                                          .readdata
			epcs_flash_controller_0_epcs_control_port_writedata  => mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_writedata,  --                                          .writedata
			epcs_flash_controller_0_epcs_control_port_chipselect => mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_chipselect, --                                          .chipselect
			green_leds_s1_address                                => mm_interconnect_0_green_leds_s1_address,                                --                             green_leds_s1.address
			green_leds_s1_write                                  => mm_interconnect_0_green_leds_s1_write,                                  --                                          .write
			green_leds_s1_readdata                               => mm_interconnect_0_green_leds_s1_readdata,                               --                                          .readdata
			green_leds_s1_writedata                              => mm_interconnect_0_green_leds_s1_writedata,                              --                                          .writedata
			green_leds_s1_chipselect                             => mm_interconnect_0_green_leds_s1_chipselect,                             --                                          .chipselect
			jtag_uart_0_avalon_jtag_slave_address                => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,                --             jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,                  --                                          .write
			jtag_uart_0_avalon_jtag_slave_read                   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,                   --                                          .read
			jtag_uart_0_avalon_jtag_slave_readdata               => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,               --                                          .readdata
			jtag_uart_0_avalon_jtag_slave_writedata              => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,              --                                          .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,            --                                          .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,             --                                          .chipselect
			key_s1_address                                       => mm_interconnect_0_key_s1_address,                                       --                                    key_s1.address
			key_s1_write                                         => mm_interconnect_0_key_s1_write,                                         --                                          .write
			key_s1_readdata                                      => mm_interconnect_0_key_s1_readdata,                                      --                                          .readdata
			key_s1_writedata                                     => mm_interconnect_0_key_s1_writedata,                                     --                                          .writedata
			key_s1_chipselect                                    => mm_interconnect_0_key_s1_chipselect,                                    --                                          .chipselect
			motor_l_s1_address                                   => mm_interconnect_0_motor_l_s1_address,                                   --                                motor_l_s1.address
			motor_l_s1_write                                     => mm_interconnect_0_motor_l_s1_write,                                     --                                          .write
			motor_l_s1_readdata                                  => mm_interconnect_0_motor_l_s1_readdata,                                  --                                          .readdata
			motor_l_s1_writedata                                 => mm_interconnect_0_motor_l_s1_writedata,                                 --                                          .writedata
			motor_l_s1_chipselect                                => mm_interconnect_0_motor_l_s1_chipselect,                                --                                          .chipselect
			motor_r_s1_address                                   => mm_interconnect_0_motor_r_s1_address,                                   --                                motor_r_s1.address
			motor_r_s1_write                                     => mm_interconnect_0_motor_r_s1_write,                                     --                                          .write
			motor_r_s1_readdata                                  => mm_interconnect_0_motor_r_s1_readdata,                                  --                                          .readdata
			motor_r_s1_writedata                                 => mm_interconnect_0_motor_r_s1_writedata,                                 --                                          .writedata
			motor_r_s1_chipselect                                => mm_interconnect_0_motor_r_s1_chipselect,                                --                                          .chipselect
			nios2_gen2_0_debug_mem_slave_address                 => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,                 --              nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                   => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,                   --                                          .write
			nios2_gen2_0_debug_mem_slave_read                    => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,                    --                                          .read
			nios2_gen2_0_debug_mem_slave_readdata                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,                --                                          .readdata
			nios2_gen2_0_debug_mem_slave_writedata               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,               --                                          .writedata
			nios2_gen2_0_debug_mem_slave_byteenable              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,              --                                          .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,             --                                          .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,             --                                          .debugaccess
			onchip_memory2_0_s1_address                          => mm_interconnect_0_onchip_memory2_0_s1_address,                          --                       onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                            => mm_interconnect_0_onchip_memory2_0_s1_write,                            --                                          .write
			onchip_memory2_0_s1_readdata                         => mm_interconnect_0_onchip_memory2_0_s1_readdata,                         --                                          .readdata
			onchip_memory2_0_s1_writedata                        => mm_interconnect_0_onchip_memory2_0_s1_writedata,                        --                                          .writedata
			onchip_memory2_0_s1_byteenable                       => mm_interconnect_0_onchip_memory2_0_s1_byteenable,                       --                                          .byteenable
			onchip_memory2_0_s1_chipselect                       => mm_interconnect_0_onchip_memory2_0_s1_chipselect,                       --                                          .chipselect
			onchip_memory2_0_s1_clken                            => mm_interconnect_0_onchip_memory2_0_s1_clken,                            --                                          .clken
			prox_sensor_s1_address                               => mm_interconnect_0_prox_sensor_s1_address,                               --                            prox_sensor_s1.address
			prox_sensor_s1_write                                 => mm_interconnect_0_prox_sensor_s1_write,                                 --                                          .write
			prox_sensor_s1_readdata                              => mm_interconnect_0_prox_sensor_s1_readdata,                              --                                          .readdata
			prox_sensor_s1_writedata                             => mm_interconnect_0_prox_sensor_s1_writedata,                             --                                          .writedata
			prox_sensor_s1_chipselect                            => mm_interconnect_0_prox_sensor_s1_chipselect,                            --                                          .chipselect
			sdram_controller_0_s1_address                        => mm_interconnect_0_sdram_controller_0_s1_address,                        --                     sdram_controller_0_s1.address
			sdram_controller_0_s1_write                          => mm_interconnect_0_sdram_controller_0_s1_write,                          --                                          .write
			sdram_controller_0_s1_read                           => mm_interconnect_0_sdram_controller_0_s1_read,                           --                                          .read
			sdram_controller_0_s1_readdata                       => mm_interconnect_0_sdram_controller_0_s1_readdata,                       --                                          .readdata
			sdram_controller_0_s1_writedata                      => mm_interconnect_0_sdram_controller_0_s1_writedata,                      --                                          .writedata
			sdram_controller_0_s1_byteenable                     => mm_interconnect_0_sdram_controller_0_s1_byteenable,                     --                                          .byteenable
			sdram_controller_0_s1_readdatavalid                  => mm_interconnect_0_sdram_controller_0_s1_readdatavalid,                  --                                          .readdatavalid
			sdram_controller_0_s1_waitrequest                    => mm_interconnect_0_sdram_controller_0_s1_waitrequest,                    --                                          .waitrequest
			sdram_controller_0_s1_chipselect                     => mm_interconnect_0_sdram_controller_0_s1_chipselect,                     --                                          .chipselect
			speaker_s1_address                                   => mm_interconnect_0_speaker_s1_address,                                   --                                speaker_s1.address
			speaker_s1_write                                     => mm_interconnect_0_speaker_s1_write,                                     --                                          .write
			speaker_s1_readdata                                  => mm_interconnect_0_speaker_s1_readdata,                                  --                                          .readdata
			speaker_s1_writedata                                 => mm_interconnect_0_speaker_s1_writedata,                                 --                                          .writedata
			speaker_s1_chipselect                                => mm_interconnect_0_speaker_s1_chipselect,                                --                                          .chipselect
			sysid_qsys_0_control_slave_address                   => mm_interconnect_0_sysid_qsys_0_control_slave_address,                   --                sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                  => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,                  --                                          .readdata
			timer_0_s1_address                                   => mm_interconnect_0_timer_0_s1_address,                                   --                                timer_0_s1.address
			timer_0_s1_write                                     => mm_interconnect_0_timer_0_s1_write,                                     --                                          .write
			timer_0_s1_readdata                                  => mm_interconnect_0_timer_0_s1_readdata,                                  --                                          .readdata
			timer_0_s1_writedata                                 => mm_interconnect_0_timer_0_s1_writedata,                                 --                                          .writedata
			timer_0_s1_chipselect                                => mm_interconnect_0_timer_0_s1_chipselect,                                --                                          .chipselect
			wifi_uart_s1_address                                 => mm_interconnect_0_wifi_uart_s1_address,                                 --                              wifi_uart_s1.address
			wifi_uart_s1_write                                   => mm_interconnect_0_wifi_uart_s1_write,                                   --                                          .write
			wifi_uart_s1_read                                    => mm_interconnect_0_wifi_uart_s1_read,                                    --                                          .read
			wifi_uart_s1_readdata                                => mm_interconnect_0_wifi_uart_s1_readdata,                                --                                          .readdata
			wifi_uart_s1_writedata                               => mm_interconnect_0_wifi_uart_s1_writedata,                               --                                          .writedata
			wifi_uart_s1_begintransfer                           => mm_interconnect_0_wifi_uart_s1_begintransfer,                           --                                          .begintransfer
			wifi_uart_s1_chipselect                              => mm_interconnect_0_wifi_uart_s1_chipselect                               --                                          .chipselect
		);

	irq_mapper : component trolley_system_irq_mapper
		port map (
			clk           => altpll_0_c0_clk,                    --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,           -- receiver5.irq
			receiver6_irq => irq_mapper_receiver6_irq,           -- receiver6.irq
			receiver7_irq => irq_mapper_receiver7_irq,           -- receiver7.irq
			sender_irq    => nios2_gen2_0_irq_irq                --    sender.irq
		);

	rst_controller : component trolley_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_001 : component trolley_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => altpll_0_c0_clk,                        --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component trolley_system_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => altpll_0_c0_clk,                    --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read_ports_inv <= not mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read;

	mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write_ports_inv <= not mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write;

	mm_interconnect_0_sdram_controller_0_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_read;

	mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_byteenable;

	mm_interconnect_0_sdram_controller_0_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_write;

	mm_interconnect_0_cam_uart_s1_read_ports_inv <= not mm_interconnect_0_cam_uart_s1_read;

	mm_interconnect_0_cam_uart_s1_write_ports_inv <= not mm_interconnect_0_cam_uart_s1_write;

	mm_interconnect_0_wifi_uart_s1_read_ports_inv <= not mm_interconnect_0_wifi_uart_s1_read;

	mm_interconnect_0_wifi_uart_s1_write_ports_inv <= not mm_interconnect_0_wifi_uart_s1_write;

	mm_interconnect_0_prox_sensor_s1_write_ports_inv <= not mm_interconnect_0_prox_sensor_s1_write;

	mm_interconnect_0_motor_r_s1_write_ports_inv <= not mm_interconnect_0_motor_r_s1_write;

	mm_interconnect_0_motor_l_s1_write_ports_inv <= not mm_interconnect_0_motor_l_s1_write;

	mm_interconnect_0_green_leds_s1_write_ports_inv <= not mm_interconnect_0_green_leds_s1_write;

	mm_interconnect_0_button_button_s1_write_ports_inv <= not mm_interconnect_0_button_button_s1_write;

	mm_interconnect_0_button_led_s1_write_ports_inv <= not mm_interconnect_0_button_led_s1_write;

	mm_interconnect_0_speaker_s1_write_ports_inv <= not mm_interconnect_0_speaker_s1_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_key_s1_write_ports_inv <= not mm_interconnect_0_key_s1_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of trolley_system
